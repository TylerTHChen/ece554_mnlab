module Bus_Interface(

);


endmodule