module tb_filter_grid();
logic clk, rst_n;



endmodule